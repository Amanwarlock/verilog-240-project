`timescale 1ns/1ns

module Bitreverse #(
	parameter DATA_WIDTH = 256
)(
	input clk,
	input enable,
	input [DATA_WIDTH-1: 0] a_in,
	output [DATA_WIDTH-1: 0] a_out
);

integer i, j;
parameter WIDTH = DATA_WIDTH-1;

reg [WIDTH: 0] res;

always @(clk or a_in or enable) begin
	if(enable === 1'b1) begin
		j = WIDTH;
		for( i = 0; i < DATA_WIDTH; i = i + 1) begin
			res[j] = a_in[i];
			j = j - 1;
		end
	
	end
end

assign a_out = res;

endmodule
